// `define NO_DELAY
`define DELAY_LEN 10
`define BUS_WIDTH 32
